module ALTERA_MF_MEMORY_INITIALIZATION;
endmodule
